parameter PIXEL_SIZE = 8;
parameter NUM_TEMPLATES = 1;
parameter LINE_SIZE = 41;
parameter NUM_OF_LINES = 34;

