parameter PIXEL_SIZE = 8;
parameter NUM_TEMPLATES = 2;
parameter LINE_SIZE = 5;
parameter NUM_OF_LINES = 5;

